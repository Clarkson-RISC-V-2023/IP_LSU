module lsu #(
    // Parameters
)(
    // Ports
);

    begin 
        // Logic definition
    end
endmodule;