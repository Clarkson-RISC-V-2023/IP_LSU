module tb_lsu #(
    // Parameters
)(
    // No_Ports
);

    begin 
        // Logic definition
    end
endmodule;